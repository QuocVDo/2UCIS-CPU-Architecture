package Definitions;
  typedef enum logic [2:0] {
    XOR,
    RXOR,
    OR,
    BEQ,
    LAND,
    MA,
    BS,
    ADDI
  } op_mne;
endpackage